library verilog;
use verilog.vl_types.all;
entity ParkingManagement_tb is
end ParkingManagement_tb;
